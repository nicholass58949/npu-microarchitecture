`include "../common/npu_definitions.vh"

module transpose_unit (
    input wire clk,
    input wire rst_n,
    
    input wire [15:0] data_in [0:63],
    input wire valid_in,
    output wire ready_in,
    output wire [15:0] data_out [0:63],
    output wire valid_out,
    input wire ready_out
);

    reg [15:0] data_out_reg [0:63];
    reg valid_out_reg;
    reg ready_in_reg;
    reg [1:0] transpose_state;

    assign data_out = data_out_reg;
    assign valid_out = valid_out_reg;
    assign ready_in = ready_in_reg;

    localparam IDLE = 2'd0;
    localparam TRANSPOSE = 2'd1;
    localparam OUTPUT = 2'd2;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (integer i = 0; i < 64; i = i + 1) begin
                data_out_reg[i] <= {16{1'b0}};
            end
            valid_out_reg <= 1'b0;
            ready_in_reg <= 1'b1;
            transpose_state <= IDLE;
        end else begin
            case (transpose_state)
                IDLE: begin
                    ready_in_reg <= 1'b1;
                    if (valid_in && ready_in_reg) begin
                        transpose_state <= TRANSPOSE;
                    end
                end
                
                TRANSPOSE: begin
                    ready_in_reg <= 1'b0;
                    for (integer i = 0; i < 8; i = i + 1) begin
                        for (integer j = 0; j < 8; j = j + 1) begin
                            data_out_reg[j * 8 + i] <= data_in[i * 8 + j];
                        end
                    end
                    transpose_state <= OUTPUT;
                end
                
                OUTPUT: begin
                    valid_out_reg <= 1'b1;
                    if (ready_out) begin
                        valid_out_reg <= 1'b0;
                        transpose_state <= IDLE;
                    end
                end
                
                default: transpose_state <= IDLE;
            endcase
        end
    end

endmodule
